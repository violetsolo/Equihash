�}�  u   ����F�Q2-(]	��� T�.!�k�~'����BϿXU�҆�1�S��Hs�hu�%{����[+�����
 MD_/U[a��>>/���g�11|/'*���ߑk����D燺�	����?繾��;�I-RY���#��F���2��/�y�'�Y˦�Z�wq�}h�z��$]��/~#I�C6�n_#��+��þG��s�������^]u�bXb��2!������J��x&^�Ǝ@4�y�7p�7�j��y(@
�H_�;j��KO���S�ә~��Pk�v,@���0��Ɠ���z=��ϝ(�\3�a�v���eX� _�z�H� =͵=Ij�s���<v%��؞t\�!#*�-!�Jܕ&>��a�q���R��g?u�����-趌)�]�'xwM��o�0�}���OIShP ��RN��$��Ro�}HɷY���UL�S��0�?H�y������FK�VH�(Fl�� ��l.b%�ڵ����#�H~߷���|�°:_UYTp�ߚ޸P����g!��u���3�	b�kf,tT�[�t�a9r��=YF�>y�A�Aq.��e������"s�B>7ʊ	�v�������mde�(�Yͭ��xA�^7^�׺W3KA�{�[+"/��F�y�����~���3j"ڼ%y��2^��;���Y�F���5�R�w8�}<K�P_��vA1cO=@�\��VO�/�\{9����i#'Fn�&RX
�(J�Itk�uL��ɭu��ɒ��̏p��R6���(��2����
�K�_��uE�@LR�D?l4�@S헱2���@��I���]r6��
^�g�>�<��-��}����=?�u�� ���K��I��6	��f0��m��Ioa���r��wA�z�]9��JUwI0|�e���l""��9���6�-�� �(�h�a�?J;���Җ��U����������62r,�F��=���:s� ���;T��l������B(
���dAB�Fj^�2��0j���Hס��ĳ[z�I^va���qH���q�jvJ�}~�4`���^`o�/�1�� �(��1��KR�8��i>3�Ճc~Pƽ3���AHm��Լ��F�y�Kw?���7`,[�Q���c�8��6x����S�~���r_�[b�%�<�|��[�L�!�[2���Sx�:�M���{�
 �*?)8���٘;�Tc:��� (���3mf�E�����[���?t<���VB�g�}��^��=	kS;vH7n�'�V�Dʉ�y��h*F��`"f�3�ˈ`�Z�X~�-a�����vX2�h��^վ������h�Ϋ?�Ff��2@�����H�>�ᣀ�1���W��,����}��1f�ZRa��ReZC�ں/q�F"K�$&84��bc�e�z�g��:�);<I���N:-˯%���U�l����a��4�"ec�(61�cJ���g�l�!�J�~p��*���7aK��G$6���0 ��m��[ؚF�����xD5|�{q���c�f�@hQ'�
�~���Z�m��A� ���Ht�/���(���jC�]�m�m�cK�����B�j�ч��=�D�d�9}�>�;��'�� �:����j=ob�m��_�[T.gP8��O/<2�7" ��3�y��p~�|i�vqu�����ng�D3��9=���YT,�N�������1���� Ϡ�Ňϲ��	f;�W����5�z������XO�īD�0��[{��	5��C:k7 �{�c��.A���H�(B�A=�g�,�M�rs@m�W$p�
3�@���Y�E�D,	�'4��	���V*�������o���D��Od~�m�^���-��\
Q�5�L�� 'N��5����|���Z�5%�)�B=e�N��ɯ��Pn��"�}�{��i�TNʈ&m��/0�JC�I�^E|<2 �]k��[�M�x��&1�slD-����q��'Tލw�n�uZ�7��F����{����duL��a]����A�Z&|�/�ic,�+/�
�F_J��C�)�	�I��I���{�&KO"�%6�ר�)��؟��P��gz.c-�rD%׈|G�K�җY�d1{���"��ƨ�U0���q�	���:d�p�8���#c�a9(���e���6��+�hF��N����%˳X�z�����K�ZL�J��M����20^��vt(IV��C�98�{䭟Ci��o{My�6-����t(JI�u�^r��IjT��Aܪ� ^�^����:��$Ê4�}~*�e�t�#��.9����7��-&v�̝5�o�}I.�V�F!}5yϼ�����Ӕ);�uc�[��@���Wk�<��� �尭�Tm��˗���u��A��b�����O#�vƿu�M�EKS�.�z�ۜwh�$VH�Iߣ��Jܻ��cyh�'޽�=�0���"�Vi5��T_��M�~�{�h�w養陲Ց�l�!�JA��r�3HP�`�R ��}��B��6������P u�=�0��MU�`�S��퓀���,�9b�UPc�lt�6���	��Q�6��(�������M?��Ɥ����
����m%�1��67.����>�;��:���
����;@e_U�Y����N=hE1��Y`GG^��bzsͨG�A!��sN�H]�BE���cq�9C���#<���t�H]]�M맮���3��c��T{�ɍ��8����bH�(��B���X*��Y���b�e��W�T��M�Q��F/��q}�>VY3��k��o��y3��B=�N�D�z
�>o,�C?M��l�:���S�!� Dx�L�_�\.�ɂH�˄^W��M��9���9�C�k9S^+����ׅ���g��9e�RV$w�W����U��`a�����?�GjЂvˌoel�N��ܤ�A��@�|d��s�^'������	��`����n�1��:�幁2��&�6���&f}�Osl�+���}�wt��W���\�Ԇ������ɿ-K&1�?�����h��WO@���g169��!ƚⲍȤ��<D�4���HBU'�-S�#Ϡ��s�!C5��A)�\
LW�
B�6���_���i!�f|����FFޱfYX*��g=c=�^]�'L����:��R���s�f+b�{�b�p}b�ܱ7{���II&^���w��jب,-u.�k�~x¥*�.�E3����*IH-�J�G�n��ΝC�W��k�A]����1t�>%�3P8)�8�����= y����r��!Z}��ȕ������AQ�6��="��_��$?>���xɩqb��1 5wC]�߈e[t�(�O�V��jar�27�k�1�S�+v&�ֈy����g��͞�P�ŜĴo8eA+�ہ�}�Lr���pa��[�̚����{t�9��҃�Î��XAQ8�AA����l�+��p1F˿b�_X�FY0��l-�K=Hm�*�+(�t@�fz�BVk�:Ț|�GЊ��kXW<�RZ���*��dԇ?bA(~ɮh�"�+�n��w�#E���虸�x!Fs�C��^���;*c}���w�JszP&���\���92���ђۦ�G�'�+��؋u_�f��8:*������M�ܮ[M�*3	��(���76�"eM~�P��3��0R���/h��73��h���J.��n�5��#�,��37l}¿�E�%��wQ�X]!�&���x2���b����Z��?�i#;-G��J�^���Q�=��N@KNR�;s�KwY�Q�C/,��R䵩�f2'�4ɤ���=�=~geX���9b٠CY�W� �� 5@�0s�����;���i�/~Ԟ�: _S��r��L���X��\�YN������RH8-;�#'�喡>:ߣ�th]��ɩ��53�^�z� ��k]]�Th"�`�3��RNjm6,�dk	���uuk8G��>E`��޵�񺟃�;l*|=L����:w|��X9
��q�����ˑVhS'c%��()�Ft
��*�aw��f\�D<�'�v�i�)n��9�o$�`Kg��m����D8ewxgUBRV�v�_��:Q�޶I����.� ��,��I=�/V�1ְ^�*���>Utw%�cb�!�\������TSd�{kfo��
�f��t%�b �1�G���gxy���,��-�	v1Zm��gBZG*"v̬x���hI��=��U�r�B�:�����KqwCvP+��;k���]���&��N+I[$��\*���T}X��e ²f�V�D�Z���-!�����M���Z	����N��}��j�t��iX=�	�δ��p�b���I6�!��UL�<L!��buR�WI��:� ^ �<3k�:�G��+
�L�S	�p�?+�H�>�S��j&Iwm�!�����e�I�S��z���
�V��ꈊ��ʿ�s�حT;�nR��0P�s��8�ه���O�$[���?�N�e&�v�� State <= S_Idle;
			end case;
		end if;
	end if;
end process;

end rtl;

