�}�  �  XHP���-(]	��� T�.!�k�~'����B/xDU�҆�1�S��H{�hu�%{����[+�����
 MD_/Ma���>/G��`�11|/+*���������o!�5(J�!=Ƞ�@�}��<���M��gMm��Q���O>a�_�GJ}�JrN~k>�Q(���l#��]b
E�Bઇ��q�Q),��妠�M(K7Fr�v[%������I�nq����S:N���:Vt3/�!x�S���D4�y�7p�7�j��y(@
�H_�;j��KO���S�ә~��Pk�v,@���0��Ɠ���z=��ϝ(�\3�a�v���eX� _�z�H� =͵=Ij�s���<v%��؞t\�!#*�-!�Jܕ&>��a�q���R��g?u�����-趌)�]�'xwM��o�0�}���OIShP ��RN��$��Ro�}HɷY���UL�S��0�?H�y������FK�VH�(Fl�� ��l�,na](t͏�詨��}@qH��R��S�Q����h"�}XQ�BnZX�%�z���^�W���'�5P��B�h����<�?�!	Ӄ>ÈF$��s�:I��P�5N^�!�n�kL�Q�/�5)��H���;�v�μB-� 8h4Ț_
'8��Y&e�d��hs� Qo	WL��>۹�]R�$��yFD @(Hhs���]MNx���w��o��Q�+GH�+$)=�!cJ!H�Z��Z���c����	�QA ��Ȟ�����c��D��p�R9�\t�峸���k ڍ��~��`�4O���#:}ho�B��ߌ�1��?ٚ��Se�������Wͨ�T�_).�Px����z�%q��"uXZ�)%g��-T 㙈��p��Jo�w����7��
��(��=��� ?�)��a=)�^���Qyw�b�j
����aMQvJ�L\Mt����Tۇ�R�\�W�Sf��M���?c��CHuINl!Jw�q�����W��R#�@ܯ��
2\�f1s�Y��$�xj��?.�U��p(���mg0L���]�ժN�\eD�p"7t,֠�[��s�AY"lm9�
j���=�'?��¯��W�"
��!�V܊��h�jMjr�?�2� ⠶[&�q��@�f� ��0�Pb�U�Z�n��A& ?$�+���٤?��Ȭ�kG>��9&U������y�J�|d��ĦF�K%=�`��e����G�nOs�����U$L�=чVb����hqY�u�N�)�Bj�m��� o	��o ��噠��x��f2���C��X�"�
&n��F�&M��j���;����p��@vO��Q��B���n�t��Y�NW۽��7� !�A%9r7-�A'_�<tR�?%�,��K���g�v�MS�?�.	�1l]�c_���Z%wB�#�D����nn���͘�-X�	��:9`*K�n�x>4ws����4�1���Ʀ�k��$�q�l�(O��}�׉X~[]������%؍�vf�9�z��n�{4�0��qĀ���x�`��]����ΟM�j_��P����'�j%�X�]��n�r�!�%ĀI�?���)���n0�MGZcMw*6��lq���������$X���P�翳��en��dy%@���άh�>���R��F���5��p>8-��HaÈ���AB���)h�]Pz�Ћ�sg��>���<��z`䑏�����Ν|w}Į�q&�Ӗ���K�Z�|maf�8"M��Q�xDGLϰ �fI�R�����r9
���M�NVdja�)*䞪��.ϵ6���o':g�
P�1��Z5����H�kd,�dyoeY._��$6u*lR?���{K\�N��Ш d@P��.A��i��:�O��s���U*>}J��3��?9�Gn��X{��:dm@g����7����]����i�����#.�z�}�ِzz.�\�#?h�7���3lD%T���>D��X�,g��;�D�A�Yɇҍ��u�2pQ��1����+s*��r�'-!��(!lS@������az�F�ʚ6�HTc- ��Yq����|�"�gvu�A���Ua%�o&o�j�l`��q	.w��hv?�YZ���;{��n��\Kʑ+.+�;Z؎��Bɐ�vL�,�hpq�f��Sn��'��M�2#��t��c�M{�H痆t�tc�Q.(��0g�j{�G�Y3�G��uÔ��"}�؇�������u��o�������8p�q^�B�(�@@�*��T5��6�xJҕ_���BS�?E��mq��]�f?�ؓn�|�\&Np[���'��R	X �ۦ�⶙��~�_�@�c�2iD�4��i����{�)(��Y�����]}��pT�=V���+����֜XRa�5�Q�%�t�1$ŋg���Yq���p�_O�`Ӣqkz��&,u�7*e�
N��3�_[�Ǧ�89�xtl�w��g!�����=�tшrValid <= '1';
					end if;
				
					
				when others => State <= S_Idle;
			end case;
		end if;
	end if;
end process;

end rtl;

