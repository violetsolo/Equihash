�}�  9   J�a����R-(]	��� T�.!�k�~'����Bϡ�_�Z�L���Gʮ[s<C�>�`�����F"���z�؁�z�O�7-Eќ����^#����LJ�Ў.��K��f�<�l1h��ߒ�Z�l$eu��]�ŗ1�U򨁼(I�t~	����mF�X5��B��x��q޴��)��M�ӟ�2)�5�����pn���H���2/�L�p�"�>�->��}��vu?.��C���{\xz�q+~d�4�y�7p�7�j��y(@
�H_�;j��KO���S�ә~��Pk�v,@���0��Ɠ���z=��ϝ(�\3�a�v���eX� _�z�H� =͵=Ij�s���<v%��؞t\�!#*�-!�Jܕ&>��a�q���R��g?u�����-趌)�]�'xwM��o�0�}���OIShP ��RN��$��Ro�}HɷY���UL�S��0�?H�y������FK�VH�(Fl�� ��l.b%��3������J~Μ�_��w�~CE�q�Q�I]}ӗٗ1�/��P�m4N�R|�G��W��;�079Nr�:��񔏃t���I6�Y�� ��=Q��O'mq�&G�_ԭ�p��ر�4����=��U�T�v�����h�8M��������{�SՁ��jh�!�#4,XǾ���%y��6l��m�ҭ$��AM� ��(�6�5rY�wa�rS��3qrS3(�;Րk[��J%���u3-K�z3*�x~�`q�MS���H�����Ш�q��v����L��(�ܸ�^�z���nL.#�YLu�:j7J�w���"�"��z��_���:B2�;�)�h�[����3������N�C��d�{��U��I�>�yeįv��e��Nle���Y��<;�I�b	
��R^OLlx�-���o"x��_���6�-�� �(�h�a�?J;���Җ��U����������62r,�F��=���:s� ���:T��l '4�Y�=~��]�L� R7Y�A�:��h�&^��)�j�-���2����:��2��׿[���r�oª
�in"ʑ������[v���J� jW���	��|�g�����GӨ�&�x�Ŕp�1T��u��*�����m~��ZS��f\O	�
�7�Q9��Cן}/��;��+oёc��Ro���X�8W����,=w� ̔�d	v�r���e��_Oq|�^� �o�e����*d��%8���M���~ځ�W$ߓʤ�"4�fS0S��x���1�Ѕ6fn\_��d�4��.���[��b��E�\�z�.��{�_�.���4;"��c��\X[+�|��cw�$/�V�I	~R�$}�(��c{�n�R��*��z��iF*���؏.�y~�w��Շ�4�4��aje����-~�;��6�n��$Dm7A��J����y6�Cڶ�kuKw,_�P�mT�_�c�y.��ܹWT{I�5C�@�|}���U�}@�Yl$R�&��j3rͰx ����yp�j�6ԣ	神ȫA�n}	�=*���K��GEB��	�(cI�j6Ԉ���k��\�ړ���>_�4�~���G���_Tl��5rqYX��B�X]���p#:�^���w���	������ ���Y�٭9�cy��3�⛊ ��DкF*�����׸�v��$� �K��&�Q�ҿ��:~���vC�o8s���Ex���/��6)�ԩ�K0�����=���]Ę��r�.D��w= �)�ni��<�i��ɀ�X^N��ٟ����t�o�ڕ���͛�+��3�'z-���X�ڽs�h,f�&�.w_�����f)�1����_L�gi�P9��ʇrN�Lm�*4A�F��6��}�V���ڱ#-j�鲯{�or�f���y$FQj�Z��X�
��޺5Fx��Wq`(�|��[`�y��8m6�����8���%�4J-ñ�/U����1LE;>�Gө������Z4�:?ʛ(�5�SlD+�sY7�Ds1��m��
�*z(�v
N�}$����"@�ʤl�È_�:��'k������}��e!����I|S�4��
֌�Bh��:L��>�'�C����\I��!�׀i�FGB��aw�G�D'�=񖴸��M���ڛL�6_�s��O �>J�G�Ta9�]�L"�!��Re>h��3��J �c@�_�o�t��t���_N��D���f�+���߰���� �2�s���8v��Yb�:�Y�,LJ�Za|D���=�m�r!w�~�.0�|���$�B|�و�Hj�vy7��z�~F��Q� ZI�-�g��Ǥt���H�C��w�r���c�k�4@�}9����:@�B<�Q[x�n,�	��!�V������(΃��9M�E>~t���{(��\�2���Û��mY�̆��tj.8�J[��ѕϑGC����"�9:����I�~3�Ol�����Z��q���`�xu���*E�4~���o�����ˢ�� (j!l�(p>=���7��@�K�RBP���O��=hXɶڼk�1��PX>�M�^�g���U=��V�d�����CF9����5z��Da��:]oK��/��H����yC��fQ��b�O	 ~[�R���#��<=G�{#i�A{C�� ��ぴ����S��Ki5���� K����KS/�����Y�_b��Rƅ��%�/�;7��j�����$vD��,[F��|w:\X,���� �n��`5�����~�ՙ`ؿ���u �{*����		��94j��#G_q$�%�"�'#�9�۠���n����]�!x"�g(����y��4ì��L�H�L7��f�T�^�QV5T��&�1uV�'�8ƫeM�l����%-������e��&7�-̺�Q���>/ۊ��o�v�����~�ky|Ž$Q6�b�>��>i��	>���士�����u�l��c�Ӛ);O��g�ݪ*���8�Ϸc��v�d�k�� )*`� 	Ӽe�l�!�J�����`Ƨ����u%m���0=���.��w���,�n2���l���H'��G�n��ܻ�jw�v�$\��*�.������ز�j����!�
����&˪&�DD�.�gN��n�D�>�;����.4�t����2_R32�l����N.gn׽xunz�imr]��|�@d�,-�a&�&l
��Բ,�Z+��U���?���gr:�OQF�vŕ������&��](ʗ���X��	.i�{���^;�^���b�e��Y0�o��~���[{��#(��P15^"��U��!Y���Pr�_�c��(�B�3~�I%��w�A�֗<�"� D�w{��Q��?���wy��|��9�ĀU�!�0aNC2�������ϡR�䁊i>�`��8�0J�W��P�\��5���S��f�-۹ó�ZV��l%Lb|�ZL�(:T�)���F��}�9bއ�v����;̢,�e��L�DslڍλFlD)�E�t��\p�O�p����`����d�H�enϲ�����2ة�dn?g;��@У|�=ΐi�YW^{aL��4�d2[z�iElIʪ:K"��edC�kH<Q<��C_Ɇ]�_�0�fg�����f%b��v���r|�#�?���Tc�K���s��U��"��	�o*-�J2����	x)��gC.��׬*���gŁ�6,���<��܏ә�bo���c�G��Rp���K3�O�^
C��~l㢰�"1�L����kF��z�X�#F����Qq��7I�o:���d�������X@������9{0�پ�3�`EK9rd2(�`��[g����q�x�n�ɒ�8S]�
JPL˹�Rĝɸ�����,�R��r� ݚ�aӐ��!��^���h{ҽ��<�jsr�z=2����"�����I�_/-�O��"@���I��������� g���<;#�r����)L?+V9ȴ	����'��@W8�S�=1(�>̏D��l#��:C���M�rհ���R�F���jgt�v��?n�.o�y�l:X�(���"p���64�n�iΈ@��������[eY��SkWtG��3�}(���P�E�N0�����`o�o��9��q�R(�8�RO��y_�{E�o�}��Us�3�_l:�uh�������TL]�f�ӭ
�s$1"����~k�;�)�NL!�<3]��4�<axH#p/w� 43��m��`����'.�Q�YICz�(T�_A�E���$t���N����Op��?_UR�6�/�,�_�9�gƟ9��>��:d��}ZV�'�K�N�5�qun��<?����sU��?�����ځq�7����X��E,��s�tq�.�n�8�blg���gIJEu��;q,��yO�nW g�i���E����Jes�yz�	�7v��-QG�)��`�n�ɦ�y�֘�h;���z
I̲�@�2ڗ���		A_�g���a
�枡Q7}ie��ue	end if;
end process;

end rtl;

