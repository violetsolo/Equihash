�}f  �   �C6[��-(]	��T�0!�k �}?W��[�vZ��e��橬�����Q
�5��S��ZL��%4U�@�_ԡw�.�Sh��A �SY�
E�>�!����'���b�E�XL}A��1�\;�寞f�Np8~Z�t%5���.0�>)��e�jt:���w��[��X(}���g�!Z�ʿl��H0����r���Mg�y���R�*�K$u��_�B�x�Y:x��\.Oxt3�D�޼���/*<���i��0M"9�2�v�5-�����B���a���q����q)ZdMT�2zv�A߼�]Y�Pk�v,@���0��Ɠ���z=��ϝ(�\3�a�v���eX� _�z�H� =͵=Ij�s���<v%��؞t\�!#*�-!�Jܕ&>��a�q���R��g?u�����-趌)�]�'xwM��o�0�}���OIShP ��RN��$��Ro�}HɷY���UL�S��0�?H�y������FK�VH�(Fl�� ��l� ��c!��i[�l(M�&x��~-�۟ՙ�tt_����k��u���\'���E8���p(M����N��X�bz�T�q��ʼ��,�D��m@wQCYH]Ӊ��A�dG�0��~e��Z3SޫZ[<v�N3�y����Y�4���k���`�^q�l1ʳS1��n�?�4�dr<b8������T]j�4��i�wp	�%�U�0V5춴d�νL��F1d�@X���� 8�rğ�į@AYٛ�P���V��Ɓ
X��Z��f/5�$jL%�"�m�PW:�}�;����ЯHj$޴8+���ŭo(��T�H$(��MgB���y4A�OK!�hVf�J�u��\`���av���_�	�(�K����E2ȀoF�+���M�)X7�H�/F:��<_4K��I4L5��͡�n���@�)���W�����$�=�̮K���&�Q�)u\\��*�F���w��M��~T�,F�M��VHu�E�!�J{�A�<�;���!N�f�өl '4�q�잨���K&�($���]�c�Tz���&��r-rrҨa�խ�9�1���;����n���L���ThʎD��S}@q]��NR�U�J&��V,�L�������Օ5��/�����C�x��u��*����60��#=�R�<�=�Pi�\e��D��.1a��YÌq&�� ���_w�ǰ2�cQ[[ǤE^��~Ji)�7ʤ�<Z/�
����9��i5 +P�W�,��f����_-��%������|�܇g#e��خ�7�Va8!�� ���%昅6fn\_��d�4��.���[��b��9��k�Z5��5�T�b�xWtz��c��\X[+�|��cw�$/�V�Iw�x,�v���+���c��7��D��Ìy�S�!â�"�(Hg	�y��H��54���p���[�b���#kvy�]KU	�1/4��T�`B���'����uCP���C��A�rs}@ΨY���D��}t��v44�݁v֬lD)�E����X0�S��kR�L%Wh���3��f>W?�����"��ŰP�-��z�����b��K��6������yӷ�^U�xڱw����H
|;�?���d~ �Bۙ���܃v��Ǐ�$�\�OJh���#Z�΀@��,G����UjOzf��t��o*-�JQ��D���;=L<��;{���Ae�ڶ�z���+���4����Ő�f��e�ޟ.̏�_5�x�j>w!��$?����{�|�η]�;8�D�g�^�3[����	l��	6S�{s��b����}���q-V������O��*G$wkR�T��S�н��U!������%IP�]	Q��-?ȗN��က��m���;�x���:D����{���'��\O扛�w�`e�m^(�'��"AF����?�SJ]f�Y�^?��gth\xn���rhk��p����B�^�_��QQ/��2g�`O͂O��-#b�c�Ao�m���Kl�%�U5���	w��N�� ��v�9���D��aMs�ϲJ��*�9NR �~����H�C��dv�+Q��%����?���N9|�����i��H�~�E�ņ9��a�w�O���x�ǯ�onf�o�{h���!4=�;h����(@;�<�c��U؊:��0�aGrd��}���X��W��	��x!In�]�'b�;b^m`��5����W�ɛ/y��aZ�|����R�G�z�hA�i��mJ�>E�l��Wnwvx|}�=i3�'��̌*�,e�f���]�_� Z��h�~��B||���W�z�H�,������ā�p��Oq��z���5\��Km�dT����EE�����..
xݯ��G�!�~pӁ,�_+�O�H�Xtw`{��So��U׈t���T�ȳ���ԐGqT�<�K���;Kȕ ���d2����'��d�W����JҷpA3Yx£=,.J�ǵ�h�\��H�m�C2=h�OȬΔ��l�,�[i0)��Y|���@}Lm�f�<��T�j�{���0<܍S�5�_H/gɭS!D�[����>��%����Xw�T�M%`�si�ڟ���)|ԩ�z�HGz��wH �O�����{�_f�j���b�ݱ���)�lwm[�#K)niБz��/�����MiT�S�P`tB�S�g���ӂ_��Ւ9���	qي��(��>G�*�����
�0�-.L���`>5������u
����,4g-�lr�~�����bk���I��j��B�[��{
���B�W�=#�c	��e��CD��AE���8e،e��;�.���-�1@#���5mg�יj����p��xƟ��p{�N�u,Mh��Bǯ	���vq�^:�̈��}n��^���~NL�U-�.V����R^�>�*�������A�{�iJ���}D��~n��+N��DM�/qY��\�R��ξ��S�1�ӵ�i��'ʻ� p"��]��X��X����9�[yl$R�&��o�c��ї�Զz(q�o�Ol�e3 Ԝ����i��%��3�ӚG�i�-�7��U.
�H�����#:e�b� +G��_p�����8E��M��S�I�Y^�)�0��L�?ɏ�q_���ɏ~���ǘ�0�c��� ���
����|_Є�zݦ����D��
T��������1���}u��4��h�B�
����h/��x;�_D�! }��9�0������V�ϿPV-��Hܸ�nY���@�����;��6a;�B� b:���
�����;������؋�b������̒�+��6�,K�m���x���f�@|�&�@!:����2	�����g�#s��q����u�?�LvT+�%l��X��|�K���܁^�݆�Un�Mrr�|3�w�]�<N�j�w0��U�¹�ל�+�&]������!��g�/�B��$_�� I�k����Y�1b�̽5E��"���!�'�(�����1n�8{'àA L��sl�$���_/O�~�3=��ɦ�8�&a0Y�M�O��>���+��)~}��d5\���&_��K��p�8�3e�_	��9%u�B-t�`�S����q���操�����~:T�F���a1 �
Nځi�f9X
<����&��~��x�~1Jz(�R�M���iB�Vh�fv߸�LaG)�Q&�3�E�\�kZ�q/ΐ����m%g�4�Uw�!CS���T<AGD7�b��%5�Փ*�t.�!six5^���!�{gN�z��<k��@��:H���Зז~�M��u6p��(*S�G,�Ƚw��;�!�N��5zf��= ���С�����FQ| ��3�1�Z�@�������n(1�Fw��:x'=QV �B�/s��T1���3�h�87�oA��$���09"�{'Nă�u�X^Y��^�1-�B8D�z��� =����h�j����p��[�Ik�(F�#=J�9q2N�b)ɇ��M!]�1�u�������&�j� �6a-�ݰ�Sl�*��Dt�H��%�-������eQ	�!J^'ɍm�͜uwT��� RL~�+m��H�Z8�*�3��9������(%(��:X]ؐ��bR��\�����ۂsf�v�AbWS,�Jd���N�K���:"�m�4| ��'�����b~�*��p�@ t�L?�V���]�!����>P���*0r�В�n���?�rC�4^l�x�D9����G�7%�1Jh����T��i\��Dׅ�g��z����΢~�p|"5����koӹ�i[MJ'ɿ�>+�&��9nkwL7\_�|z�^<�7Ɏ�,�O�NL�V�l��Kwa�#=,�WN� �aHG����զ O���U&R���@:�����ަ�����K�¼��ʸ�lɭ��![m+q
pF����$�Z�X4:Y~�5�u#��e��H��³[G�^EZ͑�&�5]��dw��.��#9����g����QS���74f���4��i�U8������ml'��a��<Υ���D.4ilO0�#�*tiz�/l��^���+��_ԥ��f�ho�]��8�q��Vd���G�X����.s�I⋢8+�և�Be("�L��!s���HI�>�a
�>q~��Z�Z�����Q�.n%ݸ̟�/��6�؎�;�'��s���,�����Zb��.|F7�r-۶ےk�n��	���Z|�Z�yc/�0�,�4�o����Os<d��&����0V�^����%��(FO6Mcߏ�z��X���C���Tյ�q(y2/�,�<��mGJz�GO�H:8㷛m�2��><o�r��͕���luЮq����-�i��>O���W��mc!z���Rz���>0�U�����v"�Q��ū��f�V�T�wG��s�Γ���&��FC-�3��+b'n��d��Y
]Ɗ�Z���5�W+�u���$� .KΪ�י\���F�ʟ�d�68������Gs�yqI�*�ğ6<Zݐ���P�E��l�$�6k4x���M�q
��*���,)E���t�S��'�c�{�W�'�N�i��tRM�`\=#-�'=�h���U�����2�B��AJ�r�r��+3-\�Ǯo
�a�P~)d��%�:4X�kNk���#W��'�I��8N%Ӆ*�k�%�ب�}$3}0�Iӄ���ʫ}��Q�������t���=g��L<X1�%k:���I�� �G��O�;)x�4R���7�`uJ�\��/��$s�R��['ᶙ���8�N����x7��Z)<
�1��^�^ �V�09�(^��WP��=�~��ۓ�E�)j,K��H]��k<<�_H����f���l!���6o`v�C���k�=��UU-9�ٓ�M�"u�x]똌�{-��n��#��Y�|�X��o��}��R�J���o|6J;1�GR��ԕ���e:.��� GQT@��@pҞ��񢱠
꺔�I���B��a@�f�����$./�zz��lD*|`�
���2�oU���Yչ�����%e�������-�"$�b=`%�ur�Y����x$+��$��؞T�"L��&=É��AK%}_s��:�:Ϥ*�^S�<�o,@�8���zL��� !�
�N�$�k9Bi�w�!�Aį�Bqx���%�!t>��߇�,p��}�5��* W32�͠�������'�/����sp^� �^+J�*sR�O�ʈ�N�&�\���1+jR
e�A�}Hҩ�������htjn⹯I5���f ���P#�y#
>1=[��gT_�my,)�p?��9��&K^�M�W%Se�
�ƛn�E^����N���1��gK�.3�M?2
�~\]�k�X�U˗NK�㾠D�% ?{b"MwT�B^ �4�j�����C��Z�Zogv�@�h�a� ��t�:LW+7N�?T��K����۩Qaw/��!|�A�Z�i=��3��Ӊ����4h�Da7����^X� {0�����T�NonWX��lD&�{����2��H�"6?�T%��_(�g���z_i<�B�2Hx��i��Ü�nʮ:�FďЊ��D
a3�p�� �kZS �YK�o���o)�R_uy>A����ڗR�Ƙ�XTJ�"q��a�^� Zlg��^6	q�(�24�d�(��J�tHg�BC�7y�q �=�z7�ȋ 9�!�l�N���hi3�����	%��7�a�<@H6W,��Ch M�y[|'�k{/����<��!�?���t#�'Hg�o��SŧI@�[y�U[y�A���J�����4�a������ؤ��N`��ClT���c0�B@Q?}�U԰V�zR������>�>k��7�fb�ڝ�{�#ꔚ����F��Y_�����C�(y*]+_y���0.�*��lԄO	_=�h���hd����j{�X����az�0���NZ��lvK��,�Vp.Ԃ����G���di��&^w�UgV�*��ω�1�bf���t]X�S)�Ţ��h�ikL~�S_mRd; -- restart read and compare process
					end if;
					
				when others => State <= S_Idle;
			end case;
		end if;
	end if;
end process;

end rtl;

