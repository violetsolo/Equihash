�}1    �d;���ԏ-(]	��� T�.��k ��'#��W��y��_"ʺEϙw�[�K��Z'ۥw�G64�����(K^��D?�I�Vk�!�#*�q�'us�ħ{��٧W�Ĉ���-�$�� .����ly�߂W�����T�6I��41�T��s8(^8k��C2]�������{��ZAX1�5zK�1�P�l�����8���*��W���!��Lۉ���wp+�Tox�Xm���({��#̀6�{�'�L�]�s��4�y�7p�7�j��y(@
�H_�;j��KO���S�ә~��Pk�v,@���0��Ɠ���z=��ϝ(�\3�a�v���eX� _�z�H� =͵=Ij�s���<v%��؞t\�!#*�-!�Jܕ&>��a�q���R��g?u�����-趌)�]�'xwM��o�0�}���OIShP ��RN��$��Ro�}HɷY���UL�S��0�?H�y������FK�VH�(Fl�� ��l�(O�����Xf[�������7����
G-B�s���50c����l�s�م�nYI±�] �0��U�
����q�R�3��|��0����>�ի��um�Up\�:����8���K8p�3z���u�	)��Zx݌�U%Y��JS
��L��a}+��#@�����=�lu`�ЗL˵���v�U�P:��b΅���h����cH�3���CN��J ^���n��LB����H�uʁiΝ+g���"r��р��k�=�6?G'�2u�T�h1�+u ��{�,�S�묌�n`ti��_�B�
* N[__�`e���ޠ9݃1毪�F:)�$H$�g���~#���!�! b�@AF,I3B��usC )l4��Fu���OQ�u���~]!,�ج5	���g��<�r�?�|]Vv�k�ƣ�5�>���ġ_K���t�~�������k�'bx��,��t��P"��#~v8�ߩd�4r9:�K����Tg��6�B�l�%�� dw�C�Z.4�ux�[�[ٝAW��T߃^|�2��d��H��A��V��V����R�q�0/���A�~ǆ��d���t.��pq�G�d�x���������~��0/����
��_R�&���gogr�0jJ�ì<+��4��Q%vZi����o{�0V!�!��ݏL�Ϧz�1�}	LщV��qi��ֽ���PT^�FOx�v=��6^4�_"�Ǐc���
�Ƅ@�9u'�?�B��b�eA7��c	���ݮl�)W�7ϓ�|���Y��m��QLJ���[ā����
_T��pd���5[�qY&���[x���@fb��G�!�}`��y����G���,��/෥B4,˪U;�k��H��di�f/UJ���'64"�����U�Ɉ0���;4.g��H��϶-��S���f���Obr:Ps�D���NC͍�5:�[��Y�*e���]��Ҡ>��$��A�=��T@�f	�by��
2�Uσ^��Q�P�Il�%�U%��!w�_����sW�!���,������l��ҹ�էv�_����Q!Ou�7�پH����'�ò���lK�MΥ�N�_��䱚TSE�4�D�H��q�.�^:� I?��3I_�/	��KlG��7*�c˦���>O��~x�ɉG�k�)>
~ܩ&��}:��v��F��Q*,Rx�T��O��=pDt4�z�c�fr������a1��O8�7�>�n�s�Rf�t��}m�m�R��Hf5r/� # .�i�rS��7�@ �I����I�i.��n�u�%��(*���C�%�2�xz���eܕ��˶w��P-W��>̉�i�Ҝ?�<��G:N�����ITͷ��L�<�~	��]�2Y�nP�..�=.<2��!�`�Fkk�:O�L��Փ�*�K���}H �`)d�k�!��b�����3G+�\�ts�M�'ySz
������@?�jm���V�S9���B�e/��mDaG8��lD+�c���s9ޑ8��\�%�;�i����/���a����w|��|��ٳc��J}�fG���X��w��q��=����v*�[���Y����T��t�����c��t�������)����R�ȆKo�ȥ�#~.L�<B+L\�yl�����)Al�آ�F0��3��m'Ò`d�3B��0��D���OR��v����B�o������ͤ�Q�^�
؄�H�%?��JP!�l�3�=]r�p3?)���V�v��!x��BW��.��$�!���!i�`6e��,�{P.��B�yS�,�Y��|�@�ȡ�s0�&��)�t�2��a�k�$@�"y���5�kR'�>O[t��\(�	��|� d��� ���l����d�KBg���i7��<X�R��	�����8���?c4�������O��j��)Qx2��T.б�{�F) �ĄN{ʀ�A��F*++��H���;{�̀��tR�w*�b�@�7�b&r���lD6-�3���S�����vTX�nT''��N��E�V.��O�U&��'���|*�(�$���*n g��7�T��=���.o@a&��Tx��jl��A�����.'��y�� n��Q7���]��PU��0��艿[�1��H��C!��9���<`4�=˕J�bށ1}*�C�	��o��#��a��^i>�aKt���ed;P�P��o�[�dp���V��Q�������Y���m�W����A;�l9P �08� �q��oiQ�`x�p}]�1s�B������>�����'���W��6{yov�Q@-�`b�Wo3?������?5���йQ �H�@��˷��%�����%+{�S����t�ZG4ҹ�}fԧ'!QBI��K��gR`I��1�`o]r�d ��g.2,DW�5�1*�$B{���`�F⅍�������4\�P<Ӓ��>&���L�]���1�������8��f,NM+���C�)�lu�j�ۺl�-	>MX@(Aݟ-��@�[�gc5�9��N�P:J����V�5�{a����#lbܞ�@{'�u{�r����M��Mo�5�:��P8)uMV�u9`:��y��2`�0�3�ୀ�8��$��f��Ub3�i:h�S)oJ Mz�)u�N��u����Yq(f^���Rg�����Kg��,�nԥƫb���7�4�',��C}����AZ��ZU�U�?q��A�t?
���u����;��*����>f�k��F�,�D"�a~*"�<�2;W4׿�݃O\��2�"�m�H���ԁ�@"%�ܮ5�ƃyw�L�l��P��=��=����^b�������
���<��5�~��N�x����&P�%iQ������ �c�|U�4 {~��B����B<r����z5)~�a���Zm�E�
٘�v��3"�`=9b�6�	�B��~���	k�U�#z��mB��/�}
X2�?C�b0aM���1���3 �t�WșZz�j��E��t�6�lD��=�>{}:������i�^P��D�s�~ͯHD�T�x!l���fꠟ�X�3�ӧe�&��4�*�j�ش۫���Z��A�i:�.A��] ����h P)�����Y���^[��l�m5m��A)��F��)������mL[� ��r�ā~�Bm�%I����*9l�d�QĪ�C�>��x҂	&p��G(]"� �Q@XUt��$��`�-��`&��f1h|~ݝ���"��<:eX#3bn7�2�m����MSʘ֡�$����e�:3�Ne�>y*:���2���������*v��$j��
3V(�m�(z�ts챿Xs�Q�K���3��h� ������.���=��Lb��^vP�6�FY��y����HwR�����p��`;2x�/k"T/\��E�9N�|!ۏ�`��P�ӻ�S�� 1�X;kO��[��F���I3"�De.��Ŗ��l�K(����~�Ó�*ud}�D�,\T�Œ��b�x5���S�{�l�&5��΀;��ۏ�#ȡF�II�����DW��;r�_d����Ҫ����p�~dJ�s2�I6�$9{���'�1k���+�O(��(�D��X_	�[�_�k��3.��7����Br[��~ܼ'��z���)�`�~H�k��.G<c�n��*Wz���5�u�*���^2��qՊr����\Q
8��;�����1E�Y��)Ҋ�b�z�2(�^���	Y݀K�P���Uq�k�\�ຕwFt�"N|�ƒTF3�)I2�P����>9���EDF���o���Y�Q��$�s��&��{\�_����հ5���~���L�w�a�̡ ��,��mCr�����rx|J��5�)(m�:E��W*�@
D�f��'^t.T@e#!������n��������G�3�	+Q�d>T~M��>��0�{��;d?��vs���ޙ�S>������s뤌�1�$�8�G��R|�ÑC��&�+�a.�b	h��y�����F�!�7l0��f&�1��-?=7v�H�����s>�tJ+)�AK���1n~�Y��s~����h�(?o��2��w�\i���N�|?�[�|�9����>�-N|�"[�9��(,e{r���<6I.67�@��tjLיM��;p1
v�tv�t"{u�wJP?��dS�O&W��Y9����,�G�XG�Q iqm��9�?t�A���v�K���ۦ~�Y��)Zڞ�,[� �ۛ��Ͼ�砿~����eS����/�Hn+����
����b��h���@5
��7t2�����	��L|����L��v��}+�b�!��t�ny�����'��n����c�"o�ڱ	
3��Ycַ��W����9������j�,rX�"`��������OG�dQn�o��n�9�1f9���'��=�,>�;��c'=2A�V��Q#���u��~~.O�`��3�>�g�:��U�^eL8���ɐ�F����)���Jg�yG�ql�(O��?C��Xf�B�y�;G��e���z���1HP��>0��k;aG��Ui`.2�UGDzI8�#��4�I.���[+zz�]��}9<��(�+��nX��l�����g�hP��/<�rZ���Ӣ����n�t}��`}O)X�f �Eh��e�<�9��D�����6�vba���F˺%���q�U�^Ut�P�~g��ܪ�?%�ɽ�C=�we#הѡg�D_G�L"!��<��[2e������t��vNMkĶ�>)��ۑ��D�a�es�}2X�6�Qo�qO# ̰4�[�T�����nB���d,uG[�)1թ��� ��Xz����-$`�JR�Y꠳h���B�E6O�Q:_��3?yLs̌;����k[�3����<LRCP�؍T-���(���#�F�2J��w�곏1�,�@]�+����T�]��x{�x��;}���L�0�~��<b����)�D]��[2y,nYn�=�4�+錵	γ_7��T�xk����l�+���M"�u��OEk�x��W�����)WY�d�6m���i*���8�����`�z--jX	o��ks�L%��%�<Nt$���栝��GN�W��t�éZ'�*�j�Ñ�O�TA�o�-�h1)`\�ׇ`��[��
�د�ٝ;,c��w�db�.PE����x�6���s�]4+�_�|�6$1�E��7v�j��Aw>R���E��yd�I{0�{�U��*�S�Y2����xD9�`�Zx��޷�%��C��?�pޢN��cv>�
gWgO�^TD�T��I�H8�	�=YS�����^"��	D1���װӭ���&x�h�ǙGk��v���"nY������lZ���HOBQk�t��tN1��k�2��k|?�wd�,��0�T�3,H2����Y����iv�ވ��V���҈o#-����Cx`y���c �Q��������%?��ZQsv"a��S��"�Ub�و��Aw��A+U�B�ZSN��d�-�0�4K7l.b%��3������H~�p��0�9�C���t/0��$(�S�2�0�^RN�w=k�Ll�m�'��9�aK9��^�v�p�]���^w���[�C�������
��0%u
���
�E�
����n�W(�]��\ؑ��Q`�b�U���Cع)̤�@:7�186 ����ƺ�%y��7\��u�����k+�y׌U��S9�r;L���l-y6=�^��mM��uzf*����s- A�g>BC�66�qZ�W@D����:�ܞ�ԳϏfā6O������%�Pţ��p�\��-.4q�
'�=i|�@?D��pk��\����|.�
�50�1O�	��9��*�C�J���(t\�q��S�m��X����pUP<��k��d��&D���+��'�.� JM��/3TO{K� ��:f^��"� ��8�h؅w��M��eH�u����	wx�T�=x۪t����m.�;���� �����e�P`��l�(O��~���Xb[uڃ-�8W�(�.�&G���g�ےIWL�\F�h���\��� ��&�MR����9�Z����w��]�\�d	��;�)>�l̶U�d^���L_.VDl�
�(��
s_��jG��f̥{f�x�
{>�q�=FJ>O@�oA�����=�db`���H��K̀�c�U�Xn��Ui�����#����h�3���p�>&�y(V��J��J?	د���I���͝b\`���sƝ�ͦ��m�4;E/�t*� �R�zE\&��l�D\������
\:S����!-e}�qW:㮀��$٘L����)*z�KS/�Q���	|����O�/,U�:49Fp�� 4B>f��&��|i8�1��ۈ=6]{T原2V���iʒY�K�m��W�X��	\��P���{Q�\�o�$#��I6�t7�N���o�GPޤ?o�������Ul��"'���f,�M��g
���4zh���&l� �\�~���n�p�Lo��#B����8�2c�\��
��b�j�ͯa�|%/)�DVz��0����ٶ�@�D �Lz��:yɞ��BN��:������|��'#�q��NM���t�T�4I�GL���=NB� =b��U���������������^���r��3�,�NJ$���#e�4��s$��J9��)����R�&@������l���עL|�Űt}KE+�B�_9�\�eb��i�ɳ�#�+dP[���e�?q`�Tz� L&��p��47rK>5�tW�\�i���Z޲l���bЕ����ݪ�^4����ܾ����q.�Z��4��@u�E<������l��W���`<E����
��B�Ty�?�a���
H��l�F����{���-!wD����,�d�<�`I�%���ju�l�+C��M�>!�6^��]����s�Fo~�V���� ��-�U�������}��t���%6f�p�`k�1Ll&��n�t��G�Y�L��>�iM�'}% ����%�aL8R:������W$��W�1�AL���oȂ�;���u�Ot�����f���3 �E%�dj�g9B�~��k�'s4\'�LZ���E@*�I�Oi���>
Z���O���ϔ���s?̤��=^(I�[���ҍ|�r�/ՉcAաk�S|�:�D� :��T��[���҂�ʏ-�c�T�m,�e0���RN�},(M]Q	��a���D�� l���"�7����_�ws�Z�&��.���؊��j�-%�Ry0�7C���;�Q���`kΤ����Fnrz�7@�&�$��Q_-ĸ�~����fa5ߑ�Mh����������3�w�^�����_r0dW�ЖMߩ�� 0 2y����]�T��1�l+Y9���6"�A�vJK�`�u�����g ��ͻk�,�9w�\M�^�Nu.�:$�6�����G�İ�t�^�c������\�a�l&����p���(�������ks
����Ý�yӗ��6I��5o �ēպ���R�N��G����.���~���T�؝������D�^��������r�r�FQ�v��u�Ѥ����]�/V���y��Ys�$��s?̤����C'	#�C���7
إM��[�tR��1"��}|-�mv�Q�{�6?\����b)���䶧��/��k�b2�w�|����D15|9����*r�o���C�]躯� �z�t�(*��z���{֎���j�%a� _�mb�[��n����/BF��̇i��ARer�x�.�~O~��G{�ø6�k����Jd&���,D��������u�V��d����\�&W^t��� )���Mv�6`%|Q,����wD����,�d�<�`I�%���ju�l�+C��M�>!�6^��]����s�Fo~�V���� ��-�U�������}��t���%6f�p�`k�1Lprocess;

end rtl;

