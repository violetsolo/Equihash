�}     @K;�X(Y-(]	��� T�.!�k�~'����B'oi4�I�d�vs���A��Y/C�>�`�����F"���z�؁�}�՛g�	��/[<�-�P���0��$	� /�}�h#g�$�`1I�ߢ�Z�l$�훷2�Nz�	�?I�D�+�DU�̷�M�pA�X5�����x�iq޴��)��-�ӟ�2Z�i1\+��%���lM(K7F���S�%������I����R��҇O��AZ���O§�p�~e�4�y�7p�7�j��y(@
�H_�;j��KO���S�ә~��Pk�v,@���0��Ɠ���z=��ϝ(�\3�a�v���eX� _�z�H� =͵=Ij�s���<v%��؞t\�!#*�-!�Jܕ&>��a�q���R��g?u�����-趌)�]�'xwM��o�0�}���OIShP ��RN��$��Ro�}HɷY���UL�S��0�?H�y������FK�VH�(Fl�� ��l�0�[{���FO����֟�0��F�7�$do�F��B����:�����^���w6�}�P�P
\
dW�Da�d:�9
�ɾ�?�~�#���1�s�	C*	���N�y��t`o�ac�^^^��l8<[����{=
L����:���Zx0��a껕���;b��V�\0Ӌ�7:�R�	h#N~�C}��4���B�ޭ��3x�pݛW���E)z� >:�w�aI�p>�bኚ%�)^!�1�nQ!+����TJ0���a��}�Kq�W��~�����P���%Y���&�/�����>S*e���^-����U"�=݄ON;�i�7}����C�Ô3tU'�{�>�	%+#���T'��=N9`/�hz����i|Ǎ9_�	sbp�D�PӛIZ��@I�Dhon��|C���6�>���n&���%���F�oB��k�ҭSO�f�e��$l�Ox�Zk7ay�������j?�U�]ie���22b�yIlD L���'�f���pau�vDc��o�}jW^� �Ԡj��V�A�=^�(cZ��$mcQ�D�h�6Ø"�=e�g �,i��Z�NyZ14	J�4x�]`_���g�hm�-�$,�ߜ�8ܭJ��W����d�EW���?���f���_���f�[��W� I��,�����p,]�E�B�v��ȟ���[ʺHyA���pᣧ5=�fH��
�>����4��O�N֟�������PF�{y�в>zˡWM�S� �%9N.�����U#��.�$����J��3��*�����Mʫ�3Zt�/-(��KoW M{�]��ur�r��[�����0��A����jӨ7�d�l����dM��l-���lD�+�1X����b�(Q��+��xB�y�(͵)�{��syh�
�\6��<��۽�خ�u�H��J���-Bh�!1�Mg	��ZKV����ѽ4)ّ6�Ew�L��ռ��k��#���*1���fc]��s��l� �\�!����WY#��[�6	�%��m&)"m�`Ͳ։c�3�ơ�rJVT*�����zc3���'����5^�q�W��ۦd�k�R;2ܑ$��H�i�H����a�q-��1����R�GL���'BX�	v��bݵ�������DW�ܜ/�����:��9�)��9� �uEi���$2�|\�����S)��M���]�?�e-���̹�6Ժ�۾J\a���
/!e�b�,�Q�w>Ԗ�죈&�bW���A�
N7�R!�P��pޏYV/&�e��sн�5�����m֏���ػR2��ɘʞ>���/�v��#d���Y'�@.I����Q8���4��`=H����Ʒ�>p5�(�(�4��]F�����d�0R�Ya���˹�mi�#]���e"g�M3��шѝ�\�����G�ޘΩ#֥��n��KЂ�@�t���큳:�R-�.y^7�F�)ݵ(��V�QI��L�8�l�%�U5���k��Y���𒜼�Y�@�w�(�@B���1<�-�� ÌG�	�?m����nJxC{g��!*J��w�+��Ҟ����sO3�;?�J��.1VvI���6Og�����(��Lco
PXǐC�oj����/�r����� ���>&7K���ͽ6j����]��rM7i�8��KG��r8M0g�l��Qq»�dێ�/m��-]�V�����m��>�S��94�$B�*��/sErnyi�y[@I�@�F1���b�x�A柳5�m�O9��h�+�y��,.�|��|M�%��.$ǹ�(���ǥ�D��$^��"Ω�(]���Qk�S`��Íj@���ú|3N:��ޢ�<�1ZL(��x�b�S�C�,9.f��-����`w�}2M�*EYv�FL���LҨ��s)�o�]D*3ahD��lXZ����Bf��ގ�8��e�w�PoTv��:?����O���`T	���dwl '4��o���t�d�.��Na'�!����h�/�x]WmA�Zxj�>W��#�����fX��[�$G?��~z���_|k �P50P��D�`�L��f�ӗj����d��:�g�Q�"�/��u��*�����rs��"+�[�/AA�Y�Bh�\$��^��.Qa����F��dܴ�[u��U�yL{��ns��<)>�XAф�yX*�;�݀�x��Z'v�0�H�F�e����I�A�Gl��δZ���}�ćk*0��ȵ�\b� /Waw��<QQ���6��5BJ7hk��8�l��.w���
��U-8���M�{�9lH�`��8�i���=g�������F=�p��sg�os\I�[�n6j �9)�v��?5�^6�f����M�9�n�ѓ*�A,%:�Э���f���WHoZ�^~Q8]�>m	�;��| ���l:����̝�ɚS�VO+�`�1r�r�͝\P�%��ј Ľ�_%���JO���jN���r Χ��a=�X�tate <= S_Wr;
						end if;
					end if;
				
				when others => State <= S_Idle;
			end case;
		end if;
	end if;
end process;

end rtl;

